-- Author: Frank Kok
-- University of Twente 2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bfar_crc_ram_B1 is
    port(
        clk				: in std_logic;
        reset			: in std_logic;
        ram_addr		: in std_logic_vector(8 downto 0); -- address to write/read ram
        ram_data_in		: in std_logic_vector(7 downto 0); -- data to write into ram
        ram_data_out	: out std_logic_vector(7 downto 0); -- data output of ram
        ram_we			: in std_logic -- write enable 
    );
    end bfar_crc_ram_B1;

architecture rtl of bfar_crc_ram_B1 is 
    type ram_array is array (511 downto 0) of std_logic_vector (7 downto 0);
signal ram: ram_array :=(
"01010000",
"00000010",
"00101111",
"00010101",
"11100000",
"10000110",
"10010101",
"11111010",
"01010001",
"00111011",
"00100100",
"10010010",
"10011111",
"00100110",
"11011000",
"00010111",
"10101110",
"11010000",
"01101100",
"11100001",
"01011001",
"10010101",
"10001111",
"00011111",
"01001100",
"01110110",
"11111001",
"00111011",
"10110110",
"00110101",
"00110001",
"01010011",
"10010001",
"01100011",
"11011110",
"00010111",
"11110111",
"01101011",
"11100110",
"01111101",
"10100000",
"10000011",
"01100011",
"10110001",
"10011001",
"00000100",
"00110110",
"10011110",
"00110010",
"10100010",
"00110001",
"01110011",
"00100100",
"10000111",
"00110100",
"10010000",
"01000010",
"00000011",
"10000100",
"01000110",
"11111010",
"01110000",
"11101100",
"01000000",
"11001000",
"01100100",
"00110110",
"10000110",
"11000001",
"00100101",
"01010011",
"00011001",
"01110110",
"10010100",
"00100011",
"10100000",
"00011101",
"00001001",
"00100010",
"01011001",
"01100000",
"00101001",
"00111001",
"11000110",
"10100000",
"11000000",
"00110010",
"00000100",
"11100011",
"11001110",
"10100000",
"00000111",
"01100000",
"10010000",
"10100110",
"10011100",
"10101111",
"11100101",
"11110111",
"01010010",
"10011010",
"00001011",
"00101000",
"00010100",
"00011011",
"00110110",
"11010100",
"01010100",
"00011111",
"01100110",
"01101010",
"10101111",
"01110101",
"00000011",
"11100001",
"01110100",
"00001010",
"01110010",
"00010100",
"00011110",
"11010101",
"10001000",
"01000000",
"11111000",
"00010000",
"11101110",
"10010001",
"00000101",
"11101100",
"00100101",
"01011010",
"11110111",
"01001100",
"01001001",
"11000010",
"01001011",
"00100000",
"10010001",
"00011000",
"10101001",
"00110111",
"01100100",
"00110101",
"00000100",
"11110011",
"01100011",
"10101000",
"00010010",
"00000000",
"00001010",
"11000100",
"01000110",
"00100010",
"11000100",
"11101001",
"00010101",
"00001111",
"00101011",
"10011111",
"11011101",
"00001001",
"01100011",
"01000000",
"10100101",
"01101011",
"01000111",
"01011001",
"11001100",
"01000011",
"10000001",
"01100100",
"00101001",
"10111000",
"10000011",
"00111000",
"01101000",
"10000000",
"11010000",
"00000111",
"11011101",
"00001000",
"00100111",
"00000010",
"11011010",
"11001001",
"00101010",
"01111001",
"00000110",
"11000111",
"10000111",
"01100110",
"01011000",
"00101011",
"00100101",
"00100111",
"01110100",
"00100001",
"10010100",
"11101010",
"10101100",
"00010010",
"10001001",
"01110111",
"10101001",
"01010001",
"00101000",
"11110101",
"10000000",
"10100010",
"10110001",
"00101001",
"01000000",
"11011100",
"00100000",
"00110010",
"10100010",
"01101100",
"10101001",
"10000010",
"10100110",
"00011111",
"11110000",
"00100100",
"01110000",
"01010000",
"10101101",
"01010100",
"10100000",
"01111000",
"10000100",
"01101101",
"10101001",
"11111100",
"11010000",
"00011101",
"11001101",
"00101011",
"00001001",
"10011011",
"01000010",
"01001110",
"00100101",
"01010110",
"00000111",
"10111010",
"11011001",
"11000000",
"11000001",
"10100000",
"01100100",
"01110111",
"10010110",
"11011101",
"11001011",
"10111000",
"00110010",
"01001100",
"01001100",
"00001111",
"10011010",
"00100010",
"00100111",
"10010010",
"00000010",
"11101100",
"11010001",
"10011000",
"01000000",
"10001110",
"10100101",
"10000101",
"11011001",
"11010010",
"00000110",
"01100101",
"11110110",
"00000010",
"01011000",
"10001001",
"10011010",
"11101100",
"01011001",
"00111010",
"10011100",
"10000010",
"01110000",
"00000110",
"01101000",
"11111101",
"11001010",
"01110000",
"11000000",
"00100010",
"10011110",
"00110000",
"00111100",
"01100101",
"10100000",
"00100000",
"10111011",
"10010001",
"00011111",
"01000100",
"10000111",
"11011011",
"01000110",
"00101011",
"10011111",
"10110011",
"00100101",
"10000010",
"10100101",
"10010011",
"01101110",
"11001001",
"01000110",
"00000010",
"01111010",
"01110000",
"11011110",
"01001001",
"10001110",
"10101100",
"11010100",
"00100110",
"10001101",
"10101100",
"11001011",
"11111010",
"10011000",
"00111010",
"10111000",
"01001000",
"00101011",
"00000001",
"01111010",
"00111100",
"10011111",
"11010001",
"00011101",
"01011110",
"10001001",
"11100010",
"00111100",
"00010101",
"01011001",
"01000001",
"10100000",
"01110000",
"11101101",
"00011101",
"10101011",
"10100010",
"00000110",
"01001000",
"00001010",
"00011100",
"00000000",
"01110000",
"10111110",
"00010101",
"10101011",
"01001010",
"01101011",
"00000111",
"00101110",
"11000100",
"00100000",
"11101100",
"00010001",
"01111011",
"10110011",
"00010101",
"11100110",
"01110001",
"00011110",
"10100100",
"00000101",
"01100010",
"10100101",
"10101101",
"10011101",
"01100001",
"00000001",
"00110111",
"01001111",
"10111011",
"10010010",
"00101011",
"00001110",
"10011000",
"11000000",
"00001000",
"00110000",
"00001101",
"11011010",
"01110110",
"11101110",
"10111000",
"00100001",
"01001010",
"10010011",
"11011110",
"00101101",
"00011101",
"01000100",
"10001001",
"11101000",
"01110111",
"10000110",
"01011101",
"01010010",
"00010011",
"11001010",
"11011010",
"00011010",
"11011001",
"10111110",
"01100110",
"11000110",
"01010001",
"11011010",
"01011001",
"01011100",
"00111001",
"00101000",
"00001010",
"00010001",
"10110111",
"11110101",
"10010111",
"01011010",
"00010100",
"00110011",
"11100111",
"10111000",
"11011101",
"10001101",
"00000111",
"00011111",
"00101010",
"01101010",
"00100010",
"00101110",
"01000001",
"01000010",
"10110100",
"11001111",
"00001010",
"00010110",
"11100100",
"10000010",
"01100000",
"10000000",
"01000110",
"10100100",
"01010010",
"00010000",
"10101001",
"01011011",
"11001100",
"00111000",
"10110100",
"00000101",
"11010101",
"00011000",
"11001010",
"10000111",
"00011001",
"10001100",
"10001000",
"11000011",
"00110010",
"00000101",
"00000001",
"01000111",
"11000110",
"01100111",
"00001000",
"01001010",
"01101001",
"01100101",
"10110010",
"00111010",
"11110000",
"11000111",
"11101110",
"11101101",
"00000011",
"10111010",
"11000110",
"01010011",
"11110001",
"01111000",
"10111001",
"01000111",
"01001010",
"10100111",
"10100100",
"01011110",
"00011101",
"11110000",
"11000011",
"01110001",
"00101000",
"11000100",
"11110100",
"01101101",
"00110011",
"00010001",
"01011101",
"01111011"
);
signal ram_out	: std_logic_vector(7 downto 0) := (others => '0');

begin 
process(clk, reset)
begin
    if rising_edge(clk) then
        if reset = '1' then
            ram_out <= (others => '0');
        else
            ram_out <= ram(to_integer(unsigned(ram_addr)));

            --Writing to ram
            if(ram_we = '1') then 
                ram(to_integer(unsigned(ram_addr))) <= ram_data_in;
            end if;
        end if;
    end if;
end process;

ram_data_out <= ram_out;

end rtl;