-- Author: Frank Kok
-- University of Twente 2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bfar_crc_ram_B0 is
    port(
        clk				: in std_logic;
        reset			: in std_logic;
        ram_addr		: in std_logic_vector(8 downto 0); -- address to write/read ram
        ram_data_in		: in std_logic_vector(7 downto 0); -- data to write into ram
        ram_data_out	: out std_logic_vector(7 downto 0); -- data output of ram
        ram_we			: in std_logic -- write enable 
    );
    end bfar_crc_ram_B0;

architecture rtl of bfar_crc_ram_B0 is 
type ram_array is array (511 downto 0) of std_logic_vector (7 downto 0);
signal ram: ram_array :=(
"01110100",
"00111000",
"01100010",
"10000100",
"10101111",
"00101010",
"01011010",
"01000000",
"10101000",
"01010000",
"11000000",
"00000001",
"00100100",
"10010111",
"10000110",
"11010100",
"10000001",
"00011011",
"00111100",
"00010010",
"00001100",
"00010001",
"11111111",
"10000011",
"10000010",
"00111001",
"00110001",
"10101100",
"11111000",
"11010011",
"00101001",
"10010100",
"10111010",
"01010101",
"10101101",
"00011010",
"00010100",
"00010101",
"00001011",
"10000110",
"00001111",
"10111001",
"00010101",
"10100010",
"00000001",
"10011000",
"11001111",
"10110001",
"10010110",
"01001100",
"00000001",
"10011100",
"00001001",
"01110000",
"00110010",
"01101000",
"00111101",
"10000111",
"01011000",
"00010001",
"10000011",
"10010100",
"01010101",
"10101000",
"01011100",
"01101111",
"11001000",
"01001011",
"00011010",
"11111111",
"01101111",
"10010111",
"00110001",
"01100100",
"00000011",
"10110100",
"10001111",
"10011100",
"00101101",
"10011000",
"00011100",
"11011000",
"10111001",
"00101001",
"10010010",
"10010111",
"10000011",
"11111000",
"11111100",
"11010111",
"11011001",
"10010011",
"10010100",
"11100101",
"00110000",
"10010000",
"10011010",
"01100000",
"11101000",
"10001100",
"00111011",
"10000100",
"11101001",
"00011001",
"01111000",
"01000001",
"10111101",
"11111001",
"00000011",
"01101001",
"00111001",
"10010100",
"00100001",
"00010001",
"10001100",
"11101011",
"00100111",
"00110000",
"00110100",
"10100011",
"00001011",
"10101101",
"01110111",
"10000111",
"11100111",
"00010100",
"10111110",
"10010001",
"10001011",
"01111010",
"00001111",
"01000000",
"10100010",
"11001100",
"11100100",
"01001011",
"01010101",
"00010001",
"01111000",
"01000110",
"00111000",
"11000011",
"00111011",
"01111010",
"00110010",
"10101101",
"11111011",
"10000111",
"01001010",
"11100001",
"10010011",
"10000010",
"01110101",
"01101001",
"11001110",
"01011011",
"10000100",
"10111101",
"10110010",
"10001110",
"01001110",
"00000011",
"10100111",
"11110101",
"01101001",
"00000000",
"10100001",
"01001001",
"11011110",
"00000011",
"01101001",
"10011001",
"00000011",
"10100000",
"00110111",
"10010110",
"11100010",
"11010011",
"11011001",
"10011110",
"00100000",
"00010000",
"11011010",
"00100001",
"00010010",
"00111000",
"01100111",
"11101100",
"11010100",
"00010011",
"10001100",
"00011010",
"01000101",
"01010000",
"00111011",
"10001010",
"11110001",
"00111111",
"10011011",
"00010010",
"11010000",
"00001110",
"00001001",
"10101010",
"10000000",
"10011100",
"01111100",
"10000100",
"11000000",
"11010011",
"11011000",
"00000001",
"10110100",
"00001101",
"11100011",
"00000100",
"11111110",
"00111101",
"00111011",
"10011110",
"00010101",
"00010001",
"01100001",
"01011000",
"01000011",
"11000000",
"00100100",
"11010110",
"00010000",
"00111010",
"10101001",
"11000110",
"00101000",
"10100100",
"01111001",
"10110011",
"00000100",
"11100100",
"10100000",
"00110001",
"11101110",
"11000001",
"11101100",
"11001001",
"00011110",
"10100000",
"10011110",
"00110000",
"10101100",
"01111000",
"01001100",
"11000111",
"10110111",
"01000000",
"11101011",
"01011001",
"10000000",
"11000000",
"11010111",
"00011010",
"00100010",
"11011010",
"10111011",
"10000100",
"11000111",
"10001001",
"00011011",
"10000100",
"10010110",
"11110001",
"10101001",
"01001101",
"00101101",
"11001000",
"01010000",
"10111000",
"01000000",
"10011110",
"11000101",
"00110111",
"10101001",
"00100010",
"11001011",
"00011110",
"01101110",
"01100010",
"11101001",
"01000100",
"11001010",
"11000000",
"00010001",
"11110001",
"00001000",
"11111001",
"10001000",
"00110010",
"00000001",
"00000010",
"11111000",
"11010011",
"10011101",
"01000001",
"00001010",
"11100100",
"00010000",
"11110000",
"11111000",
"00100010",
"10100000",
"10110110",
"10101011",
"11110110",
"10110000",
"00000001",
"00100111",
"11000101",
"00001100",
"11110111",
"11101000",
"00100010",
"00110100",
"00011101",
"00100111",
"10101001",
"00000100",
"10101101",
"11111001",
"01010100",
"10000110",
"01110000",
"11101101",
"11000001",
"11000101",
"11001001",
"00001011",
"01000101",
"10001110",
"00100010",
"00001000",
"10111001",
"00001110",
"00011100",
"01011111",
"11101111",
"10000100",
"01000101",
"01001101",
"11001110",
"01010000",
"11100011",
"10000110",
"00011110",
"10000011",
"01000000",
"00000001",
"00010010",
"11110101",
"01010010",
"11010000",
"01001010",
"00011010",
"11100100",
"00000001",
"11111110",
"10001010",
"00000000",
"10100000",
"10010000",
"11000011",
"10000100",
"01000011",
"11000100",
"11000010",
"11110001",
"10111001",
"00000010",
"11000100",
"10101001",
"11101000",
"01010010",
"10000001",
"10101111",
"01011011",
"10000000",
"00100011",
"10000101",
"00111010",
"01001111",
"01101110",
"10111001",
"10001111",
"00010011",
"10100001",
"00001100",
"10111101",
"10011100",
"01100100",
"00010011",
"10001100",
"10001011",
"10100100",
"10010011",
"11111101",
"11010011",
"10010011",
"01011100",
"00101001",
"01001110",
"11011010",
"00011011",
"10111111",
"11101101",
"11001111",
"10110001",
"11000111",
"10000100",
"01100010",
"10111101",
"10001001",
"01000011",
"00011101",
"00111100",
"00011011",
"10001101",
"10100001",
"11011111",
"00110011",
"11001000",
"11010000",
"00010010",
"01011000",
"00111010",
"11001011",
"10011111",
"10110101",
"00100001",
"00100011",
"01010000",
"10001101",
"01010000",
"01111100",
"01100111",
"11001011",
"00010001",
"00111110",
"11111000",
"01111110",
"00001101",
"10011000",
"01000100",
"00001001",
"01011011",
"01001010",
"00000011",
"00101110",
"00000000",
"10001011",
"00001001",
"10110001",
"00111011",
"10111000",
"11001101",
"01111000",
"11111110",
"10110111",
"00010010",
"01111001",
"10011110",
"11110011",
"11100001",
"01001001",
"00001010",
"01110010",
"01101001",
"01101001",
"11010110",
"10101001",
"10100001",
"00110110",
"01110100",
"00011110",
"10010001",
"00000001",
"11000000",
"11100111",
"11101001",
"00001001",
"10011000",
"10001110",
"00000111",
"11011010",
"01110000",
"00100000",
"00011100",
"10000000",
"00111100",
"10000100",
"10111010",
"10001000",
"01011000",
"01010101",
"01111111",
"00001101",
"00000001",
"01000000",
"11011110",
"01110001",
"11001100",
"01000100",
"01000000",
"00001101",
"11010111"
);
signal ram_out	: std_logic_vector(7 downto 0) := (others => '0');

begin 
process(clk, reset)
begin
    if rising_edge(clk) then
        if reset = '1' then
            ram_out <= (others => '0');
        else
            ram_out <= ram(to_integer(unsigned(ram_addr)));

            --Writing to ram
            if(ram_we = '1') then 
                ram(to_integer(unsigned(ram_addr))) <= ram_data_in;
            end if;
        end if;
    end if;
end process;

ram_data_out <= ram_out;

end rtl;