-- Author: Frank Kok
-- University of Twente 2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bfar_crc_ram_A2 is
    port(
        clk				: in std_logic;
        reset			: in std_logic;
        ram_addr		: in std_logic_vector(9 downto 0); -- address to write/read ram
        ram_data_in		: in std_logic_vector(7 downto 0); -- data to write into ram
        ram_data_out	: out std_logic_vector(7 downto 0); -- data output of ram
        ram_we			: in std_logic -- write enable 
    );
    end bfar_crc_ram_A2;

architecture rtl of bfar_crc_ram_A2 is 
type ram_array is array (1023 downto 0) of std_logic_vector (7 downto 0);
signal ram: ram_array :=(
"01111100",
"10101101",
"10111101",
"11000101",
"10000000",
"10010101",
"01100001",
"01101000",
"01000000",
"10010100",
"10011101",
"00011000",
"11011100",
"00000100",
"00010010",
"10110101",
"00010011",
"10101001",
"00001100",
"00100100",
"11000100",
"11101101",
"00000010",
"10011101",
"01100011",
"00100010",
"01001010",
"01011010",
"00110001",
"00001101",
"00001011",
"01001101",
"11001011",
"11101110",
"00001110",
"00100000",
"10110111",
"01000010",
"00101000",
"01100100",
"00110011",
"10100100",
"00101000",
"10100110",
"00110010",
"10001100",
"10110101",
"00110000",
"00010010",
"00000000",
"10000111",
"00000000",
"01010000",
"10111101",
"10001010",
"11110100",
"00010110",
"10101000",
"00000100",
"01110100",
"00101100",
"01110000",
"00010101",
"00001001",
"01000001",
"11101011",
"00000011",
"00101100",
"00000000",
"11100010",
"00001111",
"11111001",
"11100000",
"00001001",
"00000011",
"11000011",
"10100001",
"00000000",
"01010011",
"01000001",
"00000001",
"00000000",
"00111010",
"00001101",
"01000000",
"00010000",
"00001000",
"01101010",
"00110110",
"00011010",
"00000100",
"10100000",
"11000000",
"00001101",
"00101100",
"01001100",
"01101001",
"01001001",
"10110110",
"00001100",
"01011100",
"01111100",
"00000110",
"00000011",
"00000101",
"01000001",
"00111011",
"00100001",
"10001011",
"10100110",
"01000001",
"00100110",
"10110100",
"10110001",
"10010010",
"01000010",
"00010001",
"10110110",
"01010111",
"00010000",
"10101100",
"00110101",
"10010111",
"11010000",
"11110101",
"10010000",
"00100101",
"11000010",
"01001001",
"00011001",
"00110010",
"01100100",
"10011001",
"01100001",
"00100001",
"01101101",
"00001000",
"11101000",
"10100110",
"00110100",
"10001110",
"00101010",
"10000110",
"11100010",
"01100001",
"01111100",
"00001000",
"01000011",
"00000001",
"01001110",
"10111101",
"11111001",
"10000000",
"01101000",
"00000000",
"00000010",
"01001111",
"00100110",
"00100011",
"10001101",
"11010001",
"10000000",
"01000000",
"01010111",
"00011101",
"00100000",
"01000011",
"01010010",
"10101000",
"11000110",
"11001000",
"00010100",
"10111010",
"11001001",
"00011001",
"00000000",
"00101000",
"01110000",
"10100110",
"00001101",
"01101010",
"11001101",
"11000101",
"00100110",
"11000011",
"10110110",
"00110010",
"00001000",
"11100010",
"10100101",
"10000010",
"10011101",
"01001110",
"10100100",
"01010000",
"01001010",
"10100110",
"10000100",
"01010000",
"10010100",
"00000110",
"10010010",
"01000010",
"01000001",
"01010001",
"01111110",
"00010010",
"10000110",
"10001001",
"01101100",
"01000101",
"01001000",
"10100110",
"10101100",
"00000001",
"10111000",
"11000010",
"00000100",
"00000010",
"00110001",
"10000101",
"00000000",
"01011010",
"10000000",
"01110101",
"00100100",
"00011101",
"00010000",
"10000000",
"11001100",
"00001111",
"01000001",
"00000101",
"01100010",
"00001100",
"10001000",
"00000100",
"01110100",
"00110000",
"00010100",
"10111100",
"01100110",
"00001101",
"00010000",
"00101010",
"10101100",
"00011001",
"00100011",
"01000000",
"10101001",
"10010111",
"01100111",
"10101010",
"10110100",
"10010010",
"01100100",
"11000100",
"10100001",
"00000010",
"01010011",
"11110001",
"01000010",
"01010000",
"00000000",
"10001000",
"10000111",
"01101101",
"01001100",
"10001011",
"11110101",
"10010101",
"00111110",
"11010110",
"01011000",
"10001010",
"10001000",
"01000110",
"00110100",
"10000010",
"10011011",
"00000000",
"00101100",
"10110001",
"11110100",
"00110000",
"11110001",
"00000001",
"11100011",
"01000010",
"01001001",
"10010110",
"10111100",
"00111100",
"01100011",
"11001100",
"10001000",
"00000110",
"01010100",
"11000110",
"10111001",
"00101000",
"01110011",
"00011101",
"00000101",
"01111010",
"01010000",
"00001100",
"01101010",
"00100001",
"01000000",
"11010100",
"00111001",
"00000001",
"00100101",
"10000110",
"00000011",
"00001110",
"01001100",
"00110000",
"01001000",
"10000000",
"11000000",
"10001111",
"00000000",
"10100011",
"01001000",
"11010011",
"01111000",
"01010001",
"11111110",
"00001000",
"10000100",
"10000010",
"10110011",
"10010101",
"01101010",
"10000000",
"11001100",
"01000100",
"00000000",
"10110101",
"00010100",
"01001110",
"00111100",
"00001011",
"00000000",
"10010100",
"10101001",
"11001001",
"00010000",
"01001101",
"01000001",
"01001111",
"10000111",
"00101101",
"01000100",
"00100001",
"00110011",
"00001110",
"10011010",
"11111110",
"00000011",
"01000001",
"10000110",
"10001110",
"00011000",
"00001100",
"11000000",
"00100010",
"00010000",
"10001000",
"00100010",
"00110000",
"11001001",
"00100110",
"00001000",
"11101001",
"00000010",
"00001000",
"11010100",
"10100011",
"01101100",
"00101011",
"00010001",
"00000010",
"10010000",
"10001000",
"00011100",
"11011011",
"10111000",
"10001110",
"00000011",
"11010100",
"01101000",
"01000100",
"10101010",
"01001100",
"11110001",
"00110010",
"00111100",
"10010110",
"00100111",
"11100110",
"01010010",
"00010000",
"10011010",
"10101010",
"11011011",
"10110100",
"11001100",
"00000001",
"00010110",
"10011010",
"01001011",
"00000010",
"01010000",
"01001001",
"11001100",
"00100110",
"00100011",
"10011001",
"10010011",
"01001100",
"01000101",
"01101101",
"11100010",
"10101001",
"01000010",
"10001001",
"00000101",
"11000110",
"01100000",
"11110010",
"11010000",
"10110000",
"10110000",
"00001011",
"00100111",
"01011101",
"10011010",
"00010010",
"10000000",
"01100000",
"10100000",
"11011111",
"10001101",
"00000010",
"01100000",
"00010010",
"01011100",
"10100100",
"00010110",
"00000000",
"01000010",
"00110010",
"00001011",
"10010010",
"01010000",
"01000000",
"11001100",
"00111000",
"01000100",
"11000100",
"10111000",
"00100010",
"10000010",
"01000011",
"11100101",
"00111011",
"00001000",
"01000000",
"10000111",
"10100110",
"01000000",
"01011110",
"10001101",
"10000000",
"01010010",
"01110101",
"11110001",
"01100011",
"00010011",
"10101000",
"00110111",
"10100010",
"01101000",
"10011100",
"10111110",
"01101010",
"01001000",
"00000001",
"01000001",
"10000101",
"00000000",
"10100000",
"11100101",
"00010100",
"11101110",
"10011100",
"01010110",
"10100000",
"01110101",
"10000101",
"00010000",
"00010010",
"00101100",
"01011001",
"10010010",
"11100111",
"11000110",
"00101101",
"10010100",
"11101000",
"11001001",
"01101000",
"10010011",
"00001100",
"01110010",
"10001011",
"11000100",
"00100000",
"00000110",
"00111011",
"00111011",
"00111001",
"11001000",
"01000001",
"10110001",
"01001110",
"10000100",
"00101101",
"10001011",
"10101010",
"11010000",
"00100100",
"10010100",
"11000111",
"00110001",
"10100110",
"00001111",
"00100011",
"01100000",
"00000110",
"01000011",
"11000000",
"00000010",
"00011100",
"00000000",
"01010011",
"11011000",
"01010010",
"00000010",
"00000111",
"11010100",
"11000010",
"00001000",
"01000000",
"01000001",
"00000001",
"01101000",
"00001001",
"00001011",
"00101111",
"00010010",
"10110111",
"00100010",
"10001100",
"00000100",
"00110100",
"10001010",
"00000100",
"01010011",
"01100111",
"10011001",
"01011100",
"01101000",
"10001001",
"01010000",
"10100100",
"00000110",
"10001100",
"10100101",
"10110110",
"00000011",
"00001001",
"01010110",
"11000101",
"00000000",
"01110000",
"00001101",
"10100010",
"11101000",
"00101000",
"10111100",
"01001110",
"01000000",
"11101100",
"00000001",
"10101001",
"11000000",
"01010110",
"01010100",
"00101000",
"01111101",
"11101101",
"00001100",
"11000110",
"00001010",
"10101000",
"10100101",
"00101110",
"10110001",
"00000000",
"10001101",
"10000001",
"00100010",
"00111000",
"10110101",
"10111000",
"00010101",
"10011101",
"11001001",
"11100111",
"11100011",
"01110100",
"00000110",
"11110000",
"11000000",
"10001001",
"01000000",
"00011000",
"00100001",
"10000001",
"00011101",
"00100111",
"00011011",
"10000111",
"10100010",
"10010010",
"00100100",
"11100010",
"00110000",
"11010010",
"00001011",
"10011010",
"11100000",
"11001100",
"10001100",
"01101000",
"00110010",
"00101010",
"00001000",
"11110010",
"00111000",
"00000011",
"01111100",
"10100101",
"10000001",
"00100100",
"00100010",
"01000100",
"01000100",
"11100010",
"10001010",
"11011111",
"01111000",
"00000110",
"00000000",
"10010001",
"01100100",
"00010100",
"10000101",
"00100000",
"10100110",
"00011110",
"00001000",
"01110100",
"11001100",
"11100000",
"00100100",
"00010100",
"11110110",
"01010101",
"10110011",
"00101101",
"01011111",
"10010000",
"00001000",
"01010001",
"01001111",
"11000010",
"00000010",
"00001010",
"10001010",
"11110000",
"10110110",
"11110010",
"00000001",
"10100110",
"10100001",
"11000110",
"00001010",
"11001000",
"00000100",
"10100100",
"01010000",
"01101100",
"01010101",
"00110001",
"01100100",
"00100100",
"01100100",
"00011011",
"11000001",
"01101001",
"01110110",
"00100010",
"10001001",
"11100110",
"11011000",
"01010000",
"01111010",
"01100100",
"00000000",
"11010001",
"00011111",
"01010001",
"00000000",
"00100000",
"11101000",
"01011101",
"01010101",
"00111011",
"01001011",
"10011000",
"11001110",
"01000100",
"00100101",
"11110110",
"00100110",
"00101000",
"10010010",
"00001000",
"11100010",
"10010011",
"00111000",
"00000000",
"11001001",
"01100110",
"00000000",
"00010010",
"11010111",
"00011011",
"11011001",
"00001100",
"11010010",
"01100110",
"10100001",
"11110101",
"01111111",
"10100001",
"00001000",
"00000011",
"01100100",
"01000010",
"10100110",
"10000001",
"10000011",
"00011000",
"00000000",
"00110101",
"10101001",
"00011100",
"11001101",
"00100110",
"10001000",
"00111010",
"01010000",
"11101111",
"10001100",
"01000011",
"11111100",
"01000100",
"00011100",
"11100000",
"00101000",
"01000010",
"11001011",
"00010100",
"00100000",
"11000000",
"10100010",
"11110111",
"11000011",
"01100010",
"00110001",
"11100100",
"10100000",
"10001010",
"10110001",
"00111100",
"01100110",
"10000000",
"01000000",
"10001001",
"00100010",
"11101010",
"00011000",
"01010010",
"00000101",
"10100000",
"11110111",
"01011110",
"11010011",
"00101111",
"00010000",
"10110111",
"00011010",
"00010100",
"00111000",
"00001010",
"11000000",
"10001001",
"01100111",
"00110000",
"00100011",
"10100001",
"10100101",
"11001000",
"01100010",
"10111110",
"11101111",
"11010110",
"00010010",
"00110010",
"01101101",
"00100101",
"01100001",
"00010010",
"01000101",
"10000010",
"00000010",
"10000110",
"00011001",
"01011101",
"00100101",
"10100000",
"11001000",
"01111010",
"00000001",
"00001100",
"00110001",
"00101010",
"00110010",
"00100001",
"10010100",
"00000110",
"00000010",
"00000001",
"01000000",
"00001111",
"10000011",
"00001100",
"10001101",
"10001010",
"01111000",
"01000000",
"01000011",
"10100100",
"01011101",
"01001110",
"10010101",
"00000000",
"11010000",
"01011010",
"01111001",
"01001001",
"10000000",
"11101000",
"10101000",
"00111000",
"10111101",
"10100000",
"01010101",
"00011100",
"01010101",
"11000110",
"00010110",
"00111111",
"00100111",
"10000111",
"01110101",
"00010110",
"01000001",
"10010111",
"00100010",
"10010010",
"10010011",
"01011100",
"11101100",
"10000000",
"01000100",
"00000001",
"00111100",
"00010000",
"00101101",
"10000110",
"00010110",
"10100100",
"10010100",
"00110101",
"10001010",
"10000000",
"00101101",
"10110111",
"00010010",
"10010010",
"00000001",
"10010001",
"10010101",
"11000101",
"00011011",
"01000100",
"10100000",
"11100100",
"00000110",
"00101001",
"10011000",
"01000000",
"00100101",
"01000100",
"00001011",
"11101000",
"00001110",
"01000110",
"00010100",
"10000101",
"00010001",
"11000100",
"00000010",
"00100011",
"11110000",
"11001100",
"00100100",
"11011110",
"01101000",
"00000000",
"01001111",
"11110001",
"01001101",
"10000000",
"11011000",
"01000001",
"00010001",
"01110011",
"00000110",
"10101110",
"00001110",
"01100011",
"11101100",
"00110010",
"00100110",
"00000011",
"10110011",
"10001011",
"01001100",
"11100000",
"11101110",
"11001010",
"11001101",
"10000010",
"01010001",
"10000001",
"01010010",
"11110101",
"00000100",
"00000110",
"00000000",
"10101001",
"10110010",
"00100011",
"01011111",
"00010001",
"00110000",
"10010101",
"11111001",
"10010011",
"00001111",
"00000110",
"00010100",
"00101010",
"10010001",
"11010000",
"01110011",
"01011010",
"11011100",
"00111101",
"01100011",
"01000101",
"01111010",
"01011001",
"01001011",
"10110010",
"11010101",
"11010110",
"11001000",
"00111010",
"10000110",
"00110011",
"10000010",
"00010101",
"01001001",
"01111010",
"00110101",
"10000011",
"00100000",
"00011010",
"00000111",
"10000111",
"00101100",
"10001101",
"11100010",
"10100001",
"01111000"
);
signal ram_out	: std_logic_vector(7 downto 0) := (others => '0');


begin 
process(clk, reset)
begin
    if rising_edge(clk) then
        if reset = '1' then
            ram_out <= (others => '0');
        else
            ram_out <= ram(to_integer(unsigned(ram_addr)));

            --Writing to ram
            if(ram_we = '1') then 
                ram(to_integer(unsigned(ram_addr))) <= ram_data_in;
            end if;
        end if;
    end if;
end process;

ram_data_out <= ram_out;

end rtl;