-- Author: Frank Kok
-- University of Twente 2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bfar_crc_ram_A1 is
    port(
        clk				: in std_logic;
        reset			: in std_logic;
        ram_addr		: in std_logic_vector(9 downto 0); -- address to write/read ram
        ram_data_in		: in std_logic_vector(7 downto 0); -- data to write into ram
        ram_data_out	: out std_logic_vector(7 downto 0); -- data output of ram
        ram_we			: in std_logic -- write enable 
    );
    end bfar_crc_ram_A1;

architecture rtl of bfar_crc_ram_A1 is 
type ram_array is array (1023 downto 0) of std_logic_vector (7 downto 0);
signal ram: ram_array :=(
"10101000",
"00001100",
"01000000",
"00100110",
"10100000",
"11000010",
"10100001",
"00010100",
"10000001",
"00100010",
"11111010",
"11101001",
"11000100",
"10101110",
"11001100",
"00110000",
"00100001",
"00000011",
"00010001",
"01000000",
"00001011",
"00010000",
"01000010",
"00001111",
"10000100",
"10110010",
"00100100",
"10101000",
"11000111",
"00111010",
"11011101",
"00001110",
"01000101",
"00010110",
"00101010",
"10100010",
"10100100",
"00101000",
"00011001",
"00010000",
"10000111",
"00110001",
"11000110",
"10011000",
"10011000",
"00100101",
"10000010",
"00001001",
"00011100",
"00010001",
"11000000",
"11100010",
"11010111",
"10110000",
"01001001",
"00110001",
"00010101",
"01100000",
"11011000",
"10011000",
"10001100",
"00001110",
"01100011",
"00110101",
"01010110",
"10101000",
"01010000",
"00011101",
"00110100",
"10011001",
"10001010",
"11001110",
"00101001",
"11000011",
"11100000",
"01101011",
"10011110",
"00010100",
"01111000",
"01010010",
"11100001",
"00000010",
"01011100",
"10101100",
"01000000",
"10111001",
"10111111",
"00111010",
"00000000",
"11011110",
"10011110",
"10010001",
"10001101",
"11110001",
"11101100",
"00000000",
"10101000",
"10001010",
"01111000",
"00000010",
"00001101",
"10110100",
"01001000",
"10100110",
"11001001",
"00010110",
"01000000",
"00100011",
"00010001",
"10001011",
"01111000",
"01111000",
"01000111",
"11100100",
"01000001",
"01010100",
"00100110",
"11000000",
"11011000",
"00110001",
"00100001",
"01110001",
"01001001",
"10011000",
"11001010",
"00001000",
"00101010",
"00000001",
"11000010",
"01000010",
"10001000",
"10100000",
"00100100",
"00000111",
"10000101",
"01100011",
"00110110",
"00101110",
"00100111",
"00101001",
"11110000",
"01000100",
"11101101",
"01010100",
"11000101",
"00110001",
"01010111",
"10000100",
"01000001",
"01100000",
"11011110",
"00100010",
"01001011",
"01000000",
"01011101",
"00110010",
"11001000",
"11001001",
"00000010",
"10000110",
"11011111",
"00001100",
"10011011",
"00100100",
"00100010",
"00000010",
"11001100",
"11000000",
"00010100",
"10110010",
"10000011",
"01101011",
"00000101",
"00000110",
"10100111",
"00000001",
"00001100",
"10001001",
"00100000",
"10010110",
"01101000",
"00101010",
"00000101",
"01010110",
"11010010",
"01111011",
"11001011",
"01110010",
"00010011",
"01000101",
"00000010",
"00000001",
"11000111",
"01000011",
"10110110",
"11000101",
"00111110",
"11110000",
"01000000",
"01000110",
"00011110",
"10000110",
"10000000",
"01110000",
"10100000",
"10000000",
"00000000",
"10010001",
"01100101",
"00011000",
"00010001",
"10000011",
"00100000",
"01000001",
"01111100",
"10110010",
"01110011",
"00100111",
"01110011",
"00011100",
"01100011",
"10001101",
"00010000",
"10100100",
"11101100",
"01111110",
"01111001",
"00110010",
"00001011",
"01101001",
"00010011",
"11000110",
"10100000",
"00000110",
"00001010",
"11001001",
"10101100",
"10000110",
"10110110",
"01111000",
"10000110",
"10100101",
"00010010",
"10000010",
"00111000",
"00101001",
"10010110",
"11000000",
"11010011",
"01100010",
"00000110",
"00001000",
"01010110",
"00001000",
"10110100",
"10000001",
"10111000",
"01101000",
"00011101",
"00101111",
"00100110",
"10000101",
"00000100",
"01001100",
"00011111",
"10100101",
"00001000",
"11000100",
"10110100",
"01010001",
"01100000",
"01000000",
"10001110",
"10100010",
"00010011",
"10001001",
"00100010",
"00100001",
"00100001",
"11101011",
"11010010",
"01010011",
"10101100",
"00100100",
"01000001",
"01001101",
"00100110",
"01000110",
"00010110",
"00001001",
"10011011",
"10011111",
"11000011",
"01001111",
"11000100",
"00001000",
"01011010",
"10110010",
"10101000",
"00001011",
"00001011",
"10100101",
"00100010",
"01001001",
"01001010",
"10110000",
"00000010",
"10011011",
"10100010",
"11011010",
"11010111",
"00101111",
"10000110",
"10000010",
"00010000",
"00111011",
"00100100",
"00010001",
"11101110",
"00000000",
"01001101",
"00001101",
"01010010",
"00101011",
"11001101",
"00001000",
"11001011",
"01011101",
"11011110",
"10011000",
"10110110",
"01001111",
"00000000",
"10101000",
"00000011",
"10100000",
"10011000",
"00100100",
"01100001",
"01101001",
"10000010",
"11001010",
"11011000",
"00100001",
"00101110",
"11101000",
"11101010",
"11011000",
"01101010",
"10100111",
"11001110",
"00110010",
"01100000",
"10001110",
"00101110",
"00010100",
"11000111",
"00000000",
"10010011",
"01001001",
"01010010",
"10010001",
"11101000",
"01010010",
"10100000",
"11101111",
"01010101",
"00110101",
"00101000",
"11101001",
"10000011",
"11000000",
"00000010",
"00000000",
"00010011",
"00001010",
"10100110",
"01100100",
"00110001",
"00000001",
"00100111",
"01000100",
"10000100",
"10111000",
"00100010",
"00100101",
"01000000",
"00111000",
"10110000",
"00011100",
"00000110",
"00001000",
"10100110",
"00000001",
"10100100",
"10111101",
"01110000",
"01010011",
"01000001",
"11010001",
"00001000",
"10000000",
"00000111",
"00111010",
"00101010",
"11001000",
"00111010",
"10110110",
"00000001",
"11100010",
"01110110",
"01110010",
"10000010",
"11001001",
"00010010",
"01100000",
"00100001",
"10101010",
"00101011",
"01100001",
"10010101",
"10110100",
"01010011",
"11101010",
"00110000",
"11010000",
"10101000",
"01101100",
"01100011",
"01101010",
"11000101",
"10010011",
"01100010",
"00111111",
"10010101",
"10001101",
"11000010",
"10001100",
"10111000",
"01010111",
"00000111",
"00001101",
"10001100",
"01001001",
"00000100",
"10100010",
"10011010",
"11100010",
"11100100",
"10101100",
"01101000",
"00110001",
"10111110",
"01111000",
"00100010",
"01000010",
"11110000",
"00010110",
"00101100",
"10100100",
"01010101",
"10001100",
"11001100",
"01001011",
"10000010",
"00001110",
"01100011",
"00101000",
"00101100",
"00011111",
"10001000",
"10100011",
"01001000",
"10110011",
"11010010",
"01010010",
"00110000",
"10101100",
"01110111",
"00101100",
"10001110",
"10001100",
"00010000",
"10111011",
"11000010",
"01111011",
"01001001",
"10001010",
"10001100",
"01000101",
"10100010",
"00100001",
"01010000",
"01010001",
"11110010",
"01111010",
"01010000",
"11011000",
"01001001",
"11001010",
"01110101",
"01011011",
"10110001",
"01000101",
"10100001",
"00000110",
"00111000",
"00010101",
"10001010",
"11000100",
"00000000",
"00100000",
"00000100",
"00110111",
"10001110",
"00101101",
"00000001",
"10001010",
"11001100",
"01001100",
"10001100",
"00100000",
"01000100",
"01000010",
"11010000",
"00011010",
"11101011",
"00000000",
"00010100",
"01000011",
"10001110",
"10110010",
"00000001",
"10010100",
"11110000",
"01110101",
"01010011",
"01001000",
"00111010",
"00001100",
"10010101",
"10110100",
"01011010",
"11100011",
"01001011",
"11011110",
"11111101",
"01010110",
"10111001",
"11111000",
"10101100",
"00000100",
"10110110",
"01010000",
"10000110",
"00100000",
"00011110",
"10000000",
"10001000",
"10100000",
"00011100",
"01000001",
"00010101",
"01011100",
"10010100",
"01011100",
"00000111",
"01010101",
"00101001",
"00001100",
"01100011",
"00000000",
"01010101",
"10010001",
"01000010",
"11010001",
"00000110",
"00000110",
"00000101",
"01000010",
"00000010",
"00100100",
"00100000",
"01001100",
"10000011",
"00100110",
"11011000",
"01010000",
"11000101",
"01011101",
"00101011",
"00001001",
"00001101",
"11010000",
"01100011",
"01110101",
"01001101",
"00010010",
"10000000",
"11001010",
"10000110",
"10001000",
"01001010",
"00110110",
"10010001",
"00000111",
"01100010",
"10010100",
"01110010",
"00010100",
"00000111",
"11110110",
"00011000",
"11100101",
"11001101",
"00100100",
"01001110",
"10111011",
"00000000",
"00001001",
"10110000",
"00000100",
"01110011",
"11100000",
"00101111",
"10001001",
"00100110",
"11010111",
"11100001",
"00000000",
"01000000",
"01011100",
"10001110",
"10000010",
"11001001",
"10000010",
"00000111",
"10100001",
"11011000",
"00100000",
"10110011",
"00100100",
"00000000",
"11011101",
"00000111",
"10100010",
"11010100",
"11101000",
"11100110",
"11100000",
"01001100",
"01010100",
"01110100",
"00100100",
"00000101",
"10010000",
"10100101",
"00101101",
"10000001",
"10010111",
"00010011",
"11001011",
"10010010",
"10000000",
"10000001",
"10001000",
"10000010",
"01100011",
"11100000",
"10010001",
"01001101",
"01010010",
"00010010",
"00100000",
"11000001",
"01100001",
"00101110",
"10100000",
"11100100",
"10110010",
"01011101",
"00110000",
"11000011",
"10111111",
"01000101",
"00100010",
"01111101",
"00110011",
"10101001",
"00100000",
"00110010",
"10000000",
"00010001",
"00000011",
"10000110",
"10000001",
"00011011",
"01100100",
"00001001",
"10100110",
"10010100",
"01001000",
"00001000",
"11001001",
"00001011",
"01001010",
"00010100",
"00000000",
"11010001",
"00101000",
"10110010",
"01111111",
"00000101",
"11010100",
"01001001",
"01110010",
"01000011",
"00011000",
"11011110",
"11000111",
"11110000",
"00100000",
"00010100",
"11011100",
"11010000",
"00111100",
"01010001",
"10000000",
"01001110",
"00100100",
"11000100",
"10010111",
"10000001",
"10000000",
"00100101",
"10001000",
"00000001",
"01010100",
"11001000",
"11001001",
"10100001",
"01110100",
"01100101",
"00001000",
"00101100",
"11010011",
"01110010",
"10001000",
"00100000",
"10000110",
"11000100",
"10001000",
"10010110",
"01011001",
"01100011",
"00110010",
"11000001",
"00000101",
"01100000",
"01111110",
"10010001",
"01000110",
"10000010",
"00110100",
"01000110",
"01101111",
"01010001",
"01010000",
"00110100",
"10000100",
"00001011",
"10100011",
"11100001",
"10010101",
"11000000",
"01011010",
"01000010",
"00000001",
"00110001",
"10100001",
"11010000",
"10101000",
"00000110",
"01010110",
"01101010",
"01001010",
"00000000",
"00011001",
"01001110",
"01100101",
"00000100",
"00000001",
"00001100",
"00011001",
"01110000",
"11001000",
"00000010",
"11111100",
"10010011",
"00000010",
"10000011",
"10010011",
"00000000",
"01100001",
"00100011",
"01111100",
"01010110",
"01001101",
"10001110",
"01010000",
"10100100",
"10110111",
"00000101",
"11110011",
"00000110",
"00100110",
"10100100",
"00001011",
"01100000",
"00000101",
"00000000",
"00001100",
"01110001",
"11110010",
"01011010",
"01000100",
"10011110",
"10000010",
"01000010",
"00001000",
"00011001",
"00000100",
"00100011",
"00000101",
"00111000",
"00001110",
"01011000",
"00001000",
"10110011",
"11011110",
"00101100",
"00011000",
"10010110",
"10000111",
"01001011",
"01010111",
"00010010",
"00001110",
"01011001",
"11100000",
"10010001",
"01000100",
"01001100",
"01100000",
"10000001",
"11011110",
"00110110",
"10000010",
"11111010",
"00001000",
"00000001",
"11000101",
"11000000",
"00101000",
"11001001",
"00111100",
"01001100",
"10011010",
"10111100",
"00111000",
"10010000",
"10110101",
"10111100",
"00100010",
"00100001",
"00000000",
"11010010",
"00000100",
"10001001",
"10010100",
"01000010",
"00011000",
"00001011",
"10010000",
"10000000",
"00001100",
"11110001",
"00010100",
"11000100",
"00001010",
"10101010",
"11010001",
"10100100",
"11000100",
"10100100",
"01011000",
"01000000",
"01010000",
"10111111",
"00110011",
"01110101",
"11001101",
"01110010",
"00010100",
"00011010",
"00001000",
"01001101",
"11000000",
"10000110",
"00100010",
"10010011",
"10010100",
"00110000",
"01001001",
"01000100",
"00110000",
"10000011",
"01101000",
"00011000",
"10010000",
"00000010",
"00101100",
"00100010",
"01110000",
"01000101",
"00111110",
"00000000",
"01010000",
"01010010",
"01000110",
"11110001",
"00111111",
"11001000",
"00100011",
"11000000",
"10000010",
"00010011",
"11010100",
"00001000",
"10101000",
"01110001",
"11101110",
"10000001",
"10011001",
"10101101",
"01100000",
"10100000",
"11000010",
"00001111",
"10010000",
"01110111",
"11000001",
"10000001",
"00000100",
"11111010",
"11001010",
"00001110",
"10111010",
"01110011",
"01101111",
"10001011",
"01000011",
"00101100",
"00001111",
"10100111",
"00001000",
"00001101",
"11100001",
"10000000",
"00101001",
"01100100",
"10110111",
"01000000",
"01110000",
"10101100",
"11000100",
"00000011",
"00100000",
"00000110",
"00000000",
"01011011",
"00011110",
"01001100",
"01101101",
"01000011",
"00011000",
"01010110",
"01010011",
"00110000",
"11110011",
"10010101",
"10001010",
"00010000",
"10001010",
"00011001",
"01001000",
"01100000",
"00100100",
"11100000",
"00101000",
"01001001",
"00111110",
"01001100",
"01111001",
"00110110",
"01010001",
"10011000",
"00011011",
"10100001",
"10011011",
"11000100",
"01100000",
"10001000",
"01010011",
"01010111",
"01001001",
"00001000",
"00000011",
"01110000",
"11000011",
"00000100",
"01101011",
"11100000",
"11000011"
);
signal ram_out	: std_logic_vector(7 downto 0) := (others => '0');

begin 
process(clk, reset)
begin
    if rising_edge(clk) then
        if reset = '1' then
            ram_out <= (others => '0');
        else
            ram_out <= ram(to_integer(unsigned(ram_addr)));

            --Writing to ram
            if(ram_we = '1') then 
                ram(to_integer(unsigned(ram_addr))) <= ram_data_in;
            end if;
        end if;
    end if;
end process;

ram_data_out <= ram_out;

end rtl;