-- Author: Frank Kok
-- University of Twente 2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bfar_crc_ram_B2 is
    port(
        clk				: in std_logic;
        reset			: in std_logic;
        ram_addr		: in std_logic_vector(8 downto 0); -- address to write/read ram
        ram_data_in		: in std_logic_vector(7 downto 0); -- data to write into ram
        ram_data_out	: out std_logic_vector(7 downto 0); -- data output of ram
        ram_we			: in std_logic -- write enable 
    );
    end bfar_crc_ram_B2;

architecture rtl of bfar_crc_ram_B2 is 
    type ram_array is array (511 downto 0) of std_logic_vector (7 downto 0);
signal ram: ram_array :=(
"11100110",
"00100110",
"00000110",
"11001011",
"01100000",
"00011100",
"10100100",
"11111101",
"00110000",
"00111111",
"11110110",
"01111011",
"00011001",
"10011110",
"01010001",
"00011100",
"01000000",
"10001001",
"00110101",
"10101010",
"00101100",
"10001110",
"11101101",
"10110110",
"10110110",
"10100100",
"11100110",
"11000000",
"00010000",
"01010001",
"01111010",
"01010000",
"11010110",
"00011001",
"11001001",
"00111101",
"10010001",
"00000111",
"01100111",
"10001010",
"11000001",
"00111101",
"11010001",
"01111111",
"10000100",
"00001001",
"01011001",
"00111101",
"10000011",
"00100010",
"10001101",
"00001000",
"01111110",
"00010010",
"01011110",
"01001001",
"10000101",
"11010100",
"01100101",
"10101110",
"01100011",
"00000110",
"01000001",
"01000101",
"11010110",
"11100011",
"10110000",
"00100001",
"10101010",
"00110000",
"11100110",
"00011101",
"00000000",
"10010000",
"01101101",
"11000101",
"10010110",
"01001000",
"01000000",
"01010000",
"00000111",
"10001100",
"00101010",
"01111100",
"10000000",
"11001000",
"11110100",
"00011100",
"10111001",
"01101011",
"00000010",
"11010001",
"11001001",
"10100111",
"00010100",
"10100001",
"10111000",
"10111111",
"10000011",
"10101001",
"00110000",
"01111111",
"10111101",
"11011011",
"00101100",
"01100001",
"00000110",
"00001010",
"00110001",
"00000000",
"00010100",
"01011000",
"01000010",
"01011010",
"01000000",
"00000010",
"10110010",
"11001101",
"00110011",
"10010011",
"00110010",
"01010010",
"01001011",
"00001101",
"00001100",
"00011001",
"01001101",
"00010011",
"10001110",
"11100100",
"10010011",
"01000011",
"01110100",
"01000110",
"00110110",
"10111000",
"00110000",
"10000000",
"00100010",
"00110011",
"01011000",
"00001100",
"10001001",
"10100010",
"00010100",
"00000100",
"11110011",
"10000111",
"11000101",
"00111011",
"01101010",
"10001001",
"10000110",
"00111001",
"01000101",
"00100000",
"00011100",
"01110100",
"10000111",
"00101111",
"01100011",
"00000100",
"11101001",
"00101000",
"01001010",
"00010000",
"01000000",
"10100010",
"10010110",
"10101010",
"00101001",
"10000110",
"00110000",
"01101000",
"11100100",
"11111010",
"11101010",
"11100010",
"11000101",
"01111110",
"10101011",
"01101001",
"01000111",
"11100001",
"00110010",
"11101000",
"10101111",
"11000011",
"10100000",
"11110010",
"10101001",
"00000010",
"10001010",
"01101100",
"01011010",
"01110111",
"10010110",
"10100101",
"10011011",
"10010011",
"00100000",
"11000010",
"01101110",
"00111000",
"10001100",
"01001001",
"01101001",
"10100110",
"10110011",
"00011010",
"00110010",
"10010100",
"01100111",
"01010011",
"11010111",
"00111100",
"01111101",
"10110110",
"01001100",
"01100010",
"01110101",
"01100010",
"10010001",
"01100010",
"11010101",
"01001010",
"11111001",
"00111110",
"10110100",
"01010000",
"10010111",
"11011011",
"01001011",
"01111001",
"00101000",
"10101011",
"01001001",
"00000100",
"10111100",
"11000111",
"10010100",
"01101111",
"01000010",
"00110001",
"00010111",
"00111000",
"01011011",
"10011011",
"01100001",
"00010111",
"11001100",
"00000000",
"10011110",
"01001010",
"00001010",
"01110111",
"10100000",
"11100110",
"00000000",
"10110011",
"01001000",
"01110000",
"00010101",
"00000110",
"01011010",
"00001000",
"10000110",
"11011100",
"01001000",
"10011110",
"00010000",
"10111000",
"01100010",
"01111011",
"11101011",
"00101101",
"11110110",
"01111100",
"00101010",
"11101110",
"01001000",
"10011001",
"11101101",
"00110111",
"11000101",
"11011000",
"00010000",
"10000110",
"10001000",
"01001100",
"01000110",
"00111110",
"11000000",
"01101000",
"00000110",
"01101011",
"10110110",
"00010000",
"01100110",
"00101110",
"00101001",
"00101110",
"00100010",
"00010001",
"10001100",
"10000110",
"01101110",
"00111101",
"11100111",
"01111101",
"01101111",
"00011000",
"00101111",
"00110100",
"10000011",
"00101001",
"00101000",
"10001100",
"10011111",
"01011001",
"00000100",
"01110100",
"10100010",
"01010000",
"01010010",
"01010001",
"01100010",
"10001001",
"10100001",
"10100010",
"11111100",
"00100000",
"00011000",
"11110110",
"01011100",
"10010110",
"01111000",
"00000110",
"00000101",
"00100111",
"01001000",
"01100000",
"10011001",
"11001001",
"11111011",
"00011010",
"00011000",
"10010011",
"00110001",
"01110001",
"11100001",
"11111110",
"00000001",
"10110001",
"10111110",
"01101001",
"01111011",
"00110110",
"01000100",
"01101101",
"00001010",
"10001011",
"10000000",
"00100100",
"01110001",
"01110101",
"00001000",
"00010010",
"10110101",
"01001010",
"11101010",
"10011001",
"00100000",
"10010101",
"00000000",
"10110101",
"11001100",
"01101000",
"00000100",
"01010011",
"11111100",
"11111001",
"10110001",
"00011110",
"00011001",
"00011100",
"10111001",
"00101000",
"01011011",
"00011100",
"01000001",
"00010100",
"11101000",
"10000011",
"10111100",
"01110000",
"10000110",
"01001011",
"10010110",
"10101010",
"01010010",
"00001000",
"00111011",
"11011010",
"00111000",
"11110111",
"00100110",
"10111000",
"00101000",
"10001100",
"01000011",
"10010000",
"10010001",
"10000011",
"10101110",
"10110111",
"11001001",
"11101001",
"10000011",
"00100011",
"01010001",
"10111101",
"00100110",
"10000011",
"11000001",
"01011101",
"00101110",
"11000101",
"01110101",
"01111010",
"11111001",
"10011100",
"00101000",
"11010000",
"11100000",
"01011011",
"01110001",
"01000101",
"10000101",
"00001100",
"00101000",
"01011010",
"11000010",
"00001000",
"10110101",
"10101100",
"10101100",
"10111101",
"00111010",
"10000011",
"11001010",
"11000010",
"11010001",
"01101101",
"11101100",
"10111111",
"00101111",
"11110001",
"01000000",
"00001100",
"11100001",
"00100111",
"10011101",
"00001110",
"10110011",
"10010111",
"00100010",
"01100100",
"00110011",
"10101101",
"00000101",
"01000111",
"00101100",
"01010111",
"10001000",
"10101000",
"00001110",
"00111000",
"00001011",
"11101011",
"00111101",
"01010101",
"10101111",
"00100110",
"10010111",
"11110001",
"00011100",
"00111010",
"10100011",
"01010010",
"01010110",
"01111001",
"11100001",
"10011011",
"10100101",
"01111010",
"11000001",
"10000010",
"10000000",
"10000000",
"10000000",
"10100011",
"01001000",
"11010001",
"10100101",
"11010000",
"00001001",
"10010010",
"01010000",
"00100000",
"00111111",
"00101000"
);
signal ram_out	: std_logic_vector(7 downto 0) := (others => '0');

begin 
process(clk, reset)
begin
    if rising_edge(clk) then
        if reset = '1' then
            ram_out <= (others => '0');
        else
            ram_out <= ram(to_integer(unsigned(ram_addr)));

            --Writing to ram
            if(ram_we = '1') then 
                ram(to_integer(unsigned(ram_addr))) <= ram_data_in;
            end if;
        end if;
    end if;
end process;

ram_data_out <= ram_out;

end rtl;