-- Author: Frank Kok
-- University of Twente 2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bfar_crc_ram_A0 is
port(
    clk				: in std_logic;
    reset			: in std_logic;
    ram_addr		: in std_logic_vector(9 downto 0); -- address to write/read ram
    ram_data_in		: in std_logic_vector(7 downto 0); -- data to write into ram
    ram_data_out	: out std_logic_vector(7 downto 0); -- data output of ram
    ram_we			: in std_logic -- write enable 
);
end bfar_crc_ram_A0;

architecture rtl of bfar_crc_ram_A0 is 
type ram_array is array (1023 downto 0) of std_logic_vector (7 downto 0);
signal ram: ram_array :=(
"10001100",
"00000001",
"00101110",
"00000000",
"11010011",
"01000010",
"11001100",
"00010110",
"10010000",
"00000101",
"10100101",
"00010001",
"00010010",
"11001011",
"00000100",
"00001010",
"01000110",
"00110011",
"00001000",
"10110000",
"00000111",
"01000110",
"01001000",
"01001011",
"01011010",
"00111101",
"00010000",
"11000100",
"00001100",
"01011011",
"11001101",
"10000001",
"11010000",
"00111001",
"01000000",
"01100010",
"01110011",
"01010100",
"01000101",
"01101010",
"00001101",
"10100000",
"11001101",
"01010101",
"11010000",
"10001001",
"01000011",
"01111000",
"00010001",
"00010011",
"00010101",
"01001110",
"00000010",
"01001111",
"01001100",
"10000000",
"10010100",
"11000000",
"00111000",
"00100011",
"00010000",
"10011001",
"00010110",
"01101001",
"01001010",
"00101000",
"10100010",
"11001001",
"10000110",
"01000110",
"01011101",
"11010100",
"10100000",
"00101000",
"00001000",
"11110010",
"10000000",
"00000011",
"01100000",
"00101100",
"01000100",
"00110111",
"10001000",
"00110010",
"11010010",
"11001011",
"00000101",
"00000000",
"01000101",
"01110010",
"00001110",
"01000001",
"10010010",
"00010000",
"10110000",
"00100101",
"00000011",
"00000000",
"10111010",
"00010101",
"01011101",
"01000010",
"01010110",
"10000101",
"01000000",
"00000001",
"01100100",
"01000000",
"11000011",
"00010000",
"00101110",
"00111110",
"10001100",
"10010100",
"01111001",
"00111110",
"10001000",
"10100110",
"01110000",
"01000010",
"11010010",
"00010100",
"11001001",
"00100000",
"11010100",
"01110001",
"01110101",
"00000000",
"11101100",
"11111101",
"11001010",
"01001010",
"01001101",
"00101010",
"00101100",
"10001101",
"10000100",
"00111111",
"01000110",
"00001001",
"00101011",
"10000110",
"01100000",
"01001001",
"00011011",
"11010110",
"00111100",
"01100001",
"00000000",
"10001011",
"10010010",
"00000011",
"00000100",
"10010001",
"11010100",
"10010110",
"00010000",
"11000010",
"00010100",
"00010101",
"00001000",
"11110000",
"00011000",
"00001010",
"01010101",
"01111010",
"11011001",
"10100000",
"10000001",
"01000100",
"00100001",
"01010101",
"11100000",
"10000001",
"01000110",
"01000000",
"00010011",
"00011010",
"10100101",
"00101101",
"01010101",
"11110110",
"11010000",
"00101001",
"00010011",
"10010010",
"01011011",
"01000000",
"00001110",
"11011110",
"00010000",
"01001001",
"10001010",
"10001111",
"01001100",
"01000000",
"01101110",
"10010000",
"00101110",
"11111000",
"10100011",
"01011110",
"01101110",
"01111100",
"00111010",
"10010000",
"10101000",
"11000001",
"00100101",
"00010001",
"00101000",
"01100000",
"00101010",
"10011101",
"00010010",
"00101001",
"00001100",
"00011000",
"00100110",
"00111001",
"00001111",
"01000110",
"00110101",
"10010101",
"00000000",
"00011001",
"00111111",
"11001011",
"10101100",
"00001000",
"10000010",
"11011011",
"10101000",
"00111100",
"00000000",
"00110101",
"01001100",
"10011111",
"00100001",
"11110100",
"11001000",
"10101011",
"11010100",
"11101111",
"00000101",
"00011010",
"01001110",
"01000001",
"01110011",
"00100100",
"00000000",
"10111001",
"11100001",
"01110100",
"00101100",
"01000010",
"00010001",
"01010101",
"00011110",
"11001001",
"10000000",
"00010000",
"01110011",
"10001110",
"00011100",
"10000000",
"10011000",
"00011000",
"10101001",
"01110010",
"11000101",
"00010010",
"10010100",
"00010010",
"00100010",
"01111111",
"00100010",
"00011011",
"00100010",
"01000001",
"10010100",
"01011010",
"01111110",
"00010000",
"10000010",
"00000001",
"11110010",
"00011100",
"01001001",
"10011100",
"11010001",
"10010010",
"10000101",
"01001000",
"00000000",
"00100011",
"01010000",
"00100000",
"11101001",
"01101000",
"01101011",
"00000101",
"00010110",
"11000000",
"00111100",
"00010001",
"00010101",
"00011001",
"01001101",
"11100101",
"00100011",
"01010000",
"10001001",
"11000111",
"10010100",
"00110000",
"01101001",
"10010000",
"10011011",
"10001010",
"00000000",
"10111000",
"01111100",
"11000111",
"00010000",
"00001101",
"11000100",
"10010010",
"00001111",
"10000000",
"01111001",
"01000111",
"00000110",
"11011111",
"00100101",
"00000000",
"10000000",
"11000110",
"10001110",
"11010010",
"11011100",
"11001000",
"00010000",
"01111011",
"01001010",
"00010111",
"10010010",
"01011110",
"11000100",
"00101110",
"00100000",
"11000000",
"10010101",
"00001010",
"00111101",
"01000101",
"00001000",
"10110000",
"11000001",
"10101001",
"11101100",
"00010111",
"00101100",
"11111001",
"01110110",
"00000001",
"01010110",
"01010010",
"00000010",
"01010011",
"01000011",
"00010001",
"00100000",
"00110001",
"10100110",
"00001000",
"00001000",
"00011001",
"01010010",
"10111000",
"10110000",
"01000111",
"00100011",
"00000111",
"11011011",
"11111010",
"10011001",
"11000000",
"10000000",
"01101001",
"11011000",
"00001001",
"01100011",
"00000100",
"01000101",
"01010010",
"00000100",
"00010111",
"01110011",
"00001100",
"00011011",
"01001010",
"10011100",
"01011100",
"01000101",
"00000000",
"00000011",
"00000000",
"00111011",
"00110100",
"11110011",
"01100001",
"01000100",
"01111110",
"10000010",
"00110111",
"11100000",
"10100101",
"10000001",
"10111111",
"00000000",
"00010111",
"10001011",
"11010011",
"00001000",
"00001110",
"10101111",
"00101011",
"01111101",
"00100110",
"00000010",
"00000100",
"01000011",
"11100001",
"10011101",
"11001010",
"11000000",
"10011000",
"10000100",
"10000000",
"00010110",
"11101000",
"00010010",
"10100001",
"01001001",
"10110000",
"11010111",
"01100100",
"10110100",
"01000100",
"11101000",
"00001000",
"01010000",
"01010100",
"01110100",
"00000000",
"00010000",
"00100100",
"10100100",
"01010111",
"00000001",
"00000111",
"00001001",
"00101001",
"11011010",
"10100011",
"10101101",
"10101001",
"11100010",
"11111000",
"00100010",
"01101000",
"10100110",
"11110010",
"00110101",
"01110101",
"01001110",
"10000011",
"10100000",
"00101000",
"01110010",
"00000000",
"01110000",
"10010000",
"10010011",
"00110100",
"01110000",
"11110000",
"01000001",
"00011100",
"10100110",
"10110001",
"11000100",
"00100010",
"01010011",
"10101001",
"01111010",
"10000001",
"11100001",
"10111010",
"10011101",
"01001010",
"10001110",
"01110001",
"10000110",
"11010011",
"01100001",
"00000101",
"00101001",
"11010001",
"00111100",
"11100000",
"11100110",
"11101001",
"10011000",
"00010000",
"00101010",
"01011001",
"01111010",
"10000001",
"01000101",
"11011100",
"10000010",
"11100100",
"11001110",
"00000000",
"01101111",
"11001111",
"00100010",
"11101100",
"00100001",
"10110000",
"00000001",
"00011111",
"11110011",
"00000011",
"00001101",
"01011000",
"01001111",
"01010010",
"00010110",
"00100001",
"10010000",
"10001011",
"01110101",
"00100000",
"01110001",
"00001100",
"10011010",
"00101000",
"10100010",
"11001000",
"00010000",
"01011001",
"01100011",
"00000011",
"00000000",
"00010010",
"01001000",
"10110000",
"01100000",
"00100001",
"11010000",
"01100010",
"01110010",
"00000000",
"00011000",
"01010011",
"00100110",
"00011000",
"01110100",
"00011001",
"01001001",
"10111000",
"01100000",
"00001101",
"10001001",
"01111100",
"00010000",
"00110000",
"10110000",
"00000110",
"01001011",
"01010010",
"01100101",
"01000110",
"10100001",
"10001111",
"00010001",
"00011111",
"10000100",
"10011010",
"10101001",
"10010101",
"00001010",
"00001011",
"10000000",
"00111010",
"10100000",
"00010000",
"10110011",
"10000010",
"10101011",
"11000001",
"11011100",
"10111000",
"00101010",
"11000001",
"00100001",
"10100010",
"00101011",
"01000001",
"00110001",
"10101110",
"01110000",
"11100111",
"10000100",
"00111100",
"01010111",
"00100001",
"00100001",
"01010100",
"00100011",
"10000110",
"10001011",
"10110000",
"01010101",
"10000001",
"00011010",
"00010100",
"11100000",
"11100000",
"11011011",
"00010111",
"10011101",
"10010100",
"10001011",
"00000101",
"01100000",
"01000110",
"00100110",
"00110100",
"10100010",
"01100000",
"00000101",
"00000010",
"00111010",
"10000101",
"00111001",
"01110100",
"00010011",
"10001000",
"00001110",
"00001110",
"00011100",
"00000000",
"01000001",
"01111101",
"00110011",
"01010110",
"00100011",
"11011000",
"10100010",
"10101011",
"10001111",
"10010010",
"10000011",
"00001000",
"11010001",
"10000100",
"00100000",
"10110100",
"00101011",
"10101101",
"01000100",
"01001001",
"11010011",
"00000110",
"11010001",
"00000000",
"11001000",
"00100011",
"01100100",
"00011000",
"00010001",
"11011001",
"11110000",
"11000001",
"00001101",
"00100001",
"10000010",
"00000101",
"00110111",
"00111001",
"00001111",
"00000100",
"00111100",
"10000000",
"00101100",
"10110001",
"00111000",
"00010000",
"10101100",
"00101110",
"10001010",
"00111110",
"00100111",
"01010100",
"00100011",
"11001100",
"10111010",
"10000101",
"01110010",
"11010111",
"00001011",
"10010010",
"10001100",
"00000101",
"01010100",
"10001001",
"01000100",
"00000100",
"01101111",
"11100001",
"01010001",
"00100001",
"00101001",
"00010110",
"01000100",
"10100101",
"00110001",
"11100100",
"00000000",
"01101010",
"00110011",
"00100000",
"10001001",
"10000011",
"11100010",
"00010101",
"00100000",
"10110000",
"10001110",
"00111000",
"01011011",
"01110101",
"01000000",
"00100001",
"11111100",
"10101000",
"00011010",
"00101100",
"10110001",
"00001000",
"00010111",
"11000010",
"00001100",
"10001100",
"11011110",
"00000100",
"10010101",
"00010100",
"00010000",
"01110000",
"11100010",
"11100000",
"00000110",
"10001110",
"10010100",
"11010101",
"01000000",
"01101111",
"01101101",
"00000111",
"11101101",
"11010100",
"10000000",
"11011000",
"01011110",
"00011010",
"01011010",
"01101010",
"00011011",
"10000001",
"00000000",
"00100011",
"10010101",
"11010001",
"11000010",
"01000001",
"11110010",
"10100110",
"00000000",
"00000000",
"00100010",
"00000110",
"10110001",
"10010010",
"00011010",
"10011001",
"01110000",
"01011010",
"01010001",
"01100001",
"10010011",
"10010000",
"11010111",
"10010001",
"10001101",
"00111000",
"01001000",
"11010011",
"00011110",
"00000101",
"01001010",
"01011011",
"00001111",
"10001000",
"00001100",
"10110010",
"01100011",
"11010111",
"00000010",
"11001000",
"10010001",
"00000000",
"10010111",
"00011010",
"00001110",
"00110011",
"11001000",
"10001111",
"00000001",
"10100000",
"00000110",
"01001001",
"11000100",
"00110000",
"10110001",
"10100000",
"00000110",
"00100011",
"10100000",
"11001000",
"01010110",
"11000010",
"00111100",
"00110000",
"01011101",
"00111001",
"01011101",
"11111101",
"10000001",
"10000010",
"00000111",
"00001010",
"01000110",
"01100011",
"10100100",
"01100000",
"10111001",
"00010000",
"01100100",
"10110100",
"00001110",
"10011000",
"11000101",
"01100000",
"01100010",
"01101011",
"11000011",
"01001110",
"11001010",
"00100101",
"01101100",
"11111011",
"00011111",
"00010110",
"11101000",
"10001001",
"10100101",
"10100010",
"11100101",
"11100000",
"11001001",
"11000010",
"01001101",
"00010111",
"00010000",
"00001000",
"10000000",
"10001001",
"01001000",
"01001000",
"00100100",
"10001101",
"00001010",
"00000101",
"00100000",
"00100011",
"10010100",
"10111110",
"01000100",
"00101000",
"00000001",
"11000010",
"01001101",
"00000001",
"11001101",
"10001000",
"11001010",
"10110010",
"11000100",
"00010100",
"00001001",
"10001100",
"11000100",
"10000000",
"01100010",
"01001000",
"00101100",
"00010100",
"11010110",
"10001000",
"00100100",
"00010000",
"10101010",
"00001000",
"00010010",
"11100101",
"10110100",
"00000000",
"00011111",
"10010110",
"11110100",
"11100000",
"11101011",
"11010011",
"00001111",
"10000001",
"01110010",
"11111100",
"01100001",
"00001101",
"00010110",
"00001101",
"01101110",
"11001000",
"10100001",
"01011010",
"00000100",
"00010010",
"00111001",
"00001000",
"00100010",
"11110100",
"11000001",
"01101001",
"10111000",
"11010000",
"00000100",
"01000000",
"10110000",
"01100000",
"11110111",
"01001010",
"10010111",
"01100101",
"11100110",
"00010001",
"11110001",
"01100000",
"10101100",
"00011100",
"00010010",
"01110010",
"10110101",
"10101011",
"10100001",
"01110010",
"00100001",
"11010100",
"10000000",
"10100110",
"10001000",
"11111000",
"00011110",
"01111000",
"00001011",
"00100010",
"11110100",
"00001000",
"11010001",
"00011100",
"00111000",
"10100001",
"00110011",
"00000110",
"00000011",
"11101000",
"01000000",
"10100100",
"10010010",
"10000111",
"10001110",
"11001111",
"00011110",
"00100011",
"00110110",
"11000001",
"01101111",
"00000100",
"11010011",
"11101100",
"11011010",
"00100100",
"01101011",
"10101000",
"10001000",
"10001100",
"00100101",
"00111011",
"01100010",
"00011000"
);
signal ram_out	: std_logic_vector(7 downto 0) := (others => '0');

begin 
process(clk, reset)
begin
    if rising_edge(clk) then
        if reset = '1' then
            ram_out <= (others => '0');
        else
            ram_out <= ram(to_integer(unsigned(ram_addr)));

            --Writing to ram
            if(ram_we = '1') then 
                ram(to_integer(unsigned(ram_addr))) <= ram_data_in;
            end if;
        end if;
    end if;
end process;

ram_data_out <= ram_out;

end rtl;