-- Author: Frank Kok
-- University of Twente 2024
--this file contains the injected dataset that is used by the testbench

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bfar_TBmem_inj1 is
port(
    clk				: in std_logic;
    reset			: in std_logic;
    ram_addr		: in std_logic_vector(6 downto 0); -- address to write/read ram
    ram_data_in		: in std_logic_vector(63 downto 0); -- data to write into ram
    ram_data_out	: out std_logic_vector(63 downto 0); -- data output of ram
    ram_we			: in std_logic -- write enable 
);
end bfar_TBmem_inj1;

architecture rtl of bfar_TBmem_inj1 is
type ram_array is array (127 downto 0) of std_logic_vector (63 downto 0);
signal ram: ram_array :=(
    "0000000000001011000011111010000000010111100001101111011010010011",
    "0000000000001011000001111010010000000000111101101110011010110011",
    "0000000000001011000011111010101000000000100001101001011110010011",
    "0000000000001011000011111010110000000000111001101000011010110011",
    "0000000000001011000011111011000000000010110100010001111000100011",
    "0000000000001011001011111011010000000000000010101000011110010011",
    "0000000000001011000011111011100000000000000010000000011100010011",
    "0000000001001011000011111011110000000001100000010000011010010011",
    "0000000000001011001011111100000000000000110000010000011000010011",
    "0000001000001011000011111100010000000001110000010000010110010011",
    "0000000000001011000001111100100000000000000001000000010100010011",
    "0000000000001011000011111100110010101001100111111111000011111111",
    "0000000000001011000011111101000000000000000110100000101100010011",
    "0000000000001011000011111101010011110101100111111111000001101110",
    "0000000000101011000011111101100000000000010010010010100000000011",
    "0000000000001011000001111101110000000001000001110001011110010011",
    "0000000000001011000011111110000010000010101001110110010001100011",
    "0000000000001011000011111110010000000101000001110001011010010011",
    "0000000100001011000011111110100000000001000001101101011010010011",
    "0000000000001011000011111111110000000000000101101000011110010011",
    "0000000000001011000011111111000000000000100001111001011110000011",
    "0000000000001011000011111111010001010000000001111111011110010011",
    "0000000000001011000111111111100000000000100101101100011010110011",
    "0000000000001011000011111111110000000000110101111111011110110011",
    "0000000000011011000100000000000000000000110001111111011110110011",
    "0000000000001011000100000000010000000001000001101001011110010011",
    "0000000000001011000100000000100001000001000001111101010110010011",
    "0000000100001011000100000000110000000000111110000001000100100011",
    "0000000000001011000100000001000000000000000101110000111100010011",
    "0000000000001011000100000001010000000000000001011000110100010011",
    "0000000000001011000100000001100011110011010111111111010001101111",
    "0000000000001011000100000001110011111111000000010010000100010011",
    "0000000000001011000100000010000000000000001000010010000000100011",
    "0010000000001011000100000010010000000001110001010010100100000011",
    "0000000000011011000100000010100000000000100000010010010000100011",
    "0000000000001011000100000010100000000000100100010010001000100011",
    "1000000000001011000100000011000000000000000100010010011000100011",
    "0000000000001011000000000011010000000000000001010000010000010011",
    "0000000000001011000100000011100000000011000001010010110000100011",
    "0000000000001011000100000011110000000010000001011010111000100011",
    "0000000010001011000100000100000000000000000000000000010010010011",
    "0000000000001011000100000100010000000011001001001001000101100011",
    "0000000000001011000100000100100000000000110000010010000010100011",
    "0000000000001011000100000100110010000000100000010010010000000011",
    "0000000000001011000100000101000000000000010000010010011010000011",
    "0000000000001011000100000101000000000000000000010010100100000011",
    "0000000000001011000100000101100000000000000100000000010100010011",
    "0000000000001011000100000101010000000001000000010000000100010011",
    "0000000000001011000100000110000000000000000100001000000001100111",
    "0000000000001011000100000110010000000000000100000100010110010011",
    "0000000000001011000100000110100000000000100001000000010100010011",
    "0000000000001011000100000110110011000011010111111111000011101111",
    "0000000000001011000100000111000100000011100001000101010110000011",
    "0000000000001011000100000111010000001110010000100001000011101111",
    "0000000000001011001100000111100000000010101001000001110000100011",
    "0000000000001011000100000111110011111111111100100000010110010011",
    "0000000000001011000100001000000000000000000001000000010100010111",
    "0000000000001011000100001000010010111111110111110111000011101111",
    "0000000000001011000100001000100000000011100001000101010110000010",
    "0000000000001011000100001000111000001100110000000001000011101111",
    "0000000100001011000100001001000000000010101001000001110000100011",
    "0000000000001011000100001001010000000000000001001001010000100011",
    "0000100000001011000100001001100000000010101001000001110100100011",
    "0000000000001011000100001001110000000000000101011000010010010011",
    "0000000000001111000100001010000011111010010111111111000001101111",
    "0000000000000011000100001010010011111011000000010000000100010011",
    "0000000000001011000100001010100000000100100000010011010000100011",
    "0000000000001011000100001010110000000100100000010010001000100011",
    "0000000000001011000100001011000000000011001100010010111000100010",
    "0000000001001011000100001011010000000011010100010010101000100011",
    "0000000000001011000100001011100000000100100100010010011000100011",
    "0000000000001011000100001010110000000101001000010010000000100011",
    "0000000000001011000100001100000000000011010000010010110010100011",
    "0001000000001011000100001100010000000011011000010010100000100011",
    "0000000000101011000100001100100000000011011100010010011000100011",
    "0000000000001011000100001100110000000011100100010010010000100011",
    "0000000000001011000100001101000000000011100100010010001010100011",
    "0000000000001011000100001101010000000111101000010010000000100011",
    "0000000000001011000100001101100100000001101100010010111000100011",
    "0000000000001011000100001101100000000000000001010000010000010011",
    "0000010000001011000100001110000000000000000001011000100110010011",
    "0000000000001011000100001110010000000000000001101000101000010011",
    "0000000000001011000100001111100000000000000001100000010010010011",
    "0000000000001011000100101110110000000000000001100001010001100011",
    "1000000000001011000100001111000000000000000100000000010010010011",
    "0000000000001011000100001101010000000000000000000000011110010011",
    "0000000000001011000100001111100001000000000000000000100100010011",
    "0000000000001011000100001111110000100001100000000000000001101111",
    "0000000000001011000100010000010000000000000110010000100100010011",
    "0000000000001011000110010000010000000000000010010000010110010011",
    "0000000000001011000100010000110000000000000010010000010100010011",
    "0000000000001011000100010000110001100111100100000010000011111111",
    "0100000000001011000100010001000000000000001101010001011110010011",
    "0000000000001011000100010001010011111111100001111110011011100011",
    "0000000010001011000100010001100011111111111110010000100100010011",
    "0000000000001011000100010001110011111111111110011000100110011011",
    "1000000000001011000100010010000000000000000010010000010110010011",
    "0000000000001011000100010010010000000000000000010000010100010011",
    "0000000000001011000100011010100001100101110100000010000011101111",
    "0000000000001011000100010010110011111111110010011111100110010001",
    "0000000000001011000000010011000000000000000101010001101110010011",
    "0001000000001011000100010011010000000000010010011000100110010011",
    "0000001000001011000100010011100010000000000000010000110100110111",
    "0000000000001011000100010011110000000001011110011000010000010011",
    "0000000000001011000100010110000000000000000000000000110000010011",
    "0000000000001011000110010100010000000000000000000000110010010011",
    "0000000000001011000101010100100000000000000100000000101000010011",
    "0000000000001010000100010100110011111111111111010000110100010011",
    "0000000000101011000100010101000001000001011100000000011000110011",
    "0000000000001011000100011101010000001001001011001111001001100011",
    "0000000000001011000100010101100100000000000111000001101100010011",
    "0000000000001011000100010101110000000000100010010000101100110011",
    "0000000000001011000100010110100000000001001010100000110110110011",
    "0000000000001011000100010110010000000000000010100010010110010011",
    "0000000000001011000100010110100000000000000001001000010100010010",
    "0000000000001011000101010110110000000000110000010010011000100011",
    "0000000000001001000100010111000001100001010100000010000011101111",
    "0000000000001001000100010111010000000001101001010111010100110011",
    "0000000000001001000100010111100000000000110000010010011000000011",
    "0000010000001011000100010111110011111111111111110000011010110111",
    "0000100000001011000100011000000000000000000001010101100001100011",
    "0000000000001011000000011000010011111111111101010000010100010011",
    "0000000000001011000100010000100000000000110101010110010100110011",
    "0000000000001011000100011000110000000000000101010000010100010010",
    "0000000000001011010100011001000000000001000010100001011100010011",
    "0000000010001011000100011001010000000001000001110101011100010011",
    "0000000000001011000101011001100000000000101001110000011110110011",
    "0100000000001011000100011001110000000001000001111001011110010011"
);
signal ram_out	: std_logic_vector(63 downto 0) := (others => '0');

begin 
process(clk, reset)
begin
    if rising_edge(clk) then
        if reset = '1' then
            ram_out <= (others => '0');
        else
            ram_out <= ram(to_integer(unsigned(ram_addr)));

            --Writing to ram
            if(ram_we = '1') then 
                ram(to_integer(unsigned(ram_addr))) <= ram_data_in;
            end if;
        end if;
    end if;
end process;

ram_data_out <= ram_out;

end rtl;